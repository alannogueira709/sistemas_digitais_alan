library verilog;
use verilog.vl_types.all;
entity bcd_decoder_vlg_vec_tst is
end bcd_decoder_vlg_vec_tst;
